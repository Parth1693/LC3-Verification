
parameter ADD =1;
parameter AND =5;
parameter NOT =9;

parameter MODE0= 0;
parameter MODE1 =1;

parameter LD =2;
parameter LDR =6;
parameter LDI =10;

parameter LEA =14;

parameter ST =3;
parameter STR =7;
parameter STI =11;

parameter BR =0;
parameter JMP =12;